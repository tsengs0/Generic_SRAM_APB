//`include "apb_sram_config.sv"
`include "apb_sram_trans.sv"
`include "sequence/apb_sram_rw_seq.sv"
`include "sequence/apb_sram_preload_seq.sv"
`include "sequence/write_read_golden_seq.sv"
`include "apb_sram_driver.sv"
`include "apb_sram_monitor.sv"
`include "apb_sram_agent.sv"
`include "apb_sram_scoreboard.sv"
`include "apb_sram_subscriber.sv"
`include "apb_sram_env.sv"
`include "apb_sram_test.sv"